entity system is
end system;

architecture behavioral of system is
begin

end;
