entity alu is
	port(
		);
end alu;

architecture behavioral of alu is
begin
end;
